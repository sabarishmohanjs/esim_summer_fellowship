* C:\Users\sabarishmohan\eSim-Workspace\54f64_test\54f64_test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/09/25 12:13:51

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U2-Pad1_ Net-_U4-Pad10_ Net-_U4-Pad9_ Net-_U4-Pad8_ Net-_U4-Pad7_ Net-_U4-Pad6_ ic_54f64		
U4  B0 C0 D0 A3 B3 Net-_U4-Pad6_ Net-_U4-Pad7_ Net-_U4-Pad8_ Net-_U4-Pad9_ Net-_U4-Pad10_ adc_bridge_5		
U1  A0 A2 B2 A1 B1 C1 Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ adc_bridge_6		
U2  Net-_U2-Pad1_ out dac_bridge_1		
R1  out GND 1k		
U3  out plot_v1		
v11  B0 GND pulse		
v10  C0 GND pulse		
v9  D0 GND pulse		
v8  A3 GND pulse		
v7  B3 GND pulse		
v6  C1 GND pulse		
v5  B1 GND pulse		
v4  A1 GND pulse		
v3  B2 GND pulse		
v2  A2 GND pulse		
v1  A0 GND pulse		
U5  A0 plot_v1		
U6  A2 plot_v1		
U7  B2 plot_v1		
U8  A1 plot_v1		
U9  B1 plot_v1		
U11  B3 plot_v1		
U12  A3 plot_v1		
U13  D0 plot_v1		
U14  C0 plot_v1		
U15  B0 plot_v1		
U10  C1 plot_v1		

.end
