* C:\FOSSEE\eSim\library\SubcircuitLibrary\54f64\54f64.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/22/25 13:59:39

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U6  Net-_U1-Pad3_ Net-_U1-Pad2_ Net-_U2-Pad1_ d_and		
X1  Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U2-Pad2_ 3_and		
U5  Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U4-Pad1_ d_and		
U4  Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U3-Pad1_ d_nor		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ d_nor		
U3  Net-_U3-Pad1_ Net-_U2-Pad3_ Net-_U1-Pad8_ d_nor		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ PORT		
X2  Net-_U1-Pad13_ Net-_U1-Pad12_ Net-_U1-Pad11_ Net-_U1-Pad1_ Net-_U4-Pad2_ 4_and		

.end
