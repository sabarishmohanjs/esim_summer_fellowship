* C:\FOSSEE\eSim\library\SubcircuitLibrary\cd4077b\cd4077b.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/24/25 14:56:23

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M3  Net-_M11-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad1_ Net-_M11-Pad1_ eSim_MOS_P		
M2  Net-_M2-Pad1_ Net-_M2-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M4  Net-_M11-Pad1_ Net-_M2-Pad2_ Net-_M2-Pad1_ Net-_M11-Pad1_ eSim_MOS_P		
M6  Net-_M1-Pad1_ Net-_M2-Pad1_ Net-_M10-Pad2_ Net-_M11-Pad1_ eSim_MOS_P		
M5  Net-_M1-Pad1_ Net-_M2-Pad2_ Net-_M10-Pad2_ Net-_M1-Pad3_ eSim_MOS_N		
M7  Net-_M10-Pad2_ Net-_M1-Pad1_ Net-_M7-Pad3_ Net-_M7-Pad3_ eSim_MOS_N		
M9  Net-_M2-Pad1_ Net-_M1-Pad1_ Net-_M10-Pad2_ Net-_M11-Pad1_ eSim_MOS_P		
M8  Net-_M7-Pad3_ Net-_M2-Pad1_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M10  Net-_M10-Pad1_ Net-_M10-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M11  Net-_M11-Pad1_ Net-_M10-Pad2_ Net-_M10-Pad1_ Net-_M11-Pad1_ eSim_MOS_P		
U1  Net-_M2-Pad2_ Net-_M1-Pad2_ Net-_M10-Pad1_ Net-_M10-Pad1_ Net-_M1-Pad2_ Net-_M2-Pad2_ Net-_M1-Pad3_ Net-_M2-Pad2_ Net-_M1-Pad2_ Net-_M10-Pad1_ Net-_M10-Pad1_ Net-_M1-Pad2_ Net-_M2-Pad2_ Net-_M11-Pad1_ PORT		

.end
